module and_3_tb();
reg a,b,c;
wire d;
and_3_gate DUT(a,b,c,d);
initial
    begin
    a=0;b=0;c=0;
    #10;
    a=0;b=0;c=1;
    #10;
    a=0;b=1;c=0;
    #10;
    a=0;b=1;c=1;
    #10;
    a=1;b=0;c=0;
    #10;
    a=1;b=0;c=1;
    #10;
    a=1;b=1;c=0;
    #10;
    a=1;b=1;c=1;
    #10;
    $finish(1);
    end
initial
    begin
    $dumpfile("test.vcd");
    $dumpvars(1);
    end
initial
    begin
    $monitor("a=%b b=%b c=%b d=%b",a,b,c,d);
    end
endmodule
