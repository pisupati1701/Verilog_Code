module and_3_gate(input wire a,b,c,output wire d);
assign temp=a&b;
assign d=temp&c;
endmodule
